module cv32e40s_miter (
  input clk,
  input rst,
  output logic alert_major_o_1,
  output logic alert_major_o_2,
  output logic alert_minor_o_1,
  output logic alert_minor_o_2,
  input logic[31:0] boot_addr_i_1,
  input logic[31:0] boot_addr_i_2,
  input logic clic_irq_i_1,
  input logic clic_irq_i_2,
  input logic[4:0] clic_irq_id_i_1,
  input logic[4:0] clic_irq_id_i_2,
  input logic[7:0] clic_irq_level_i_1,
  input logic[7:0] clic_irq_level_i_2,
  input logic[1:0] clic_irq_priv_i_1,
  input logic[1:0] clic_irq_priv_i_2,
  input logic clic_irq_shv_i_1,
  input logic clic_irq_shv_i_2,
  output logic core_sleep_o_1,
  output logic core_sleep_o_2,
  output logic[12:0] data_achk_o_1,
  output logic[12:0] data_achk_o_2,
  output logic[31:0] data_addr_o_1,
  output logic[31:0] data_addr_o_2,
  output logic[3:0] data_be_o_1,
  output logic[3:0] data_be_o_2,
  output logic data_dbg_o_1,
  output logic data_dbg_o_2,
  input logic data_err_i_1,
  input logic data_err_i_2,
  input logic data_gnt_i_1,
  input logic data_gnt_i_2,
  input logic data_gntpar_i_1,
  input logic data_gntpar_i_2,
  output logic[1:0] data_memtype_o_1,
  output logic[1:0] data_memtype_o_2,
  output logic[2:0] data_prot_o_1,
  output logic[2:0] data_prot_o_2,
  input logic[4:0] data_rchk_i_1,
  input logic[4:0] data_rchk_i_2,
  input logic[31:0] data_rdata_i_1,
  input logic[31:0] data_rdata_i_2,
  output logic data_req_o_1,
  output logic data_req_o_2,
  output logic data_reqpar_o_1,
  output logic data_reqpar_o_2,
  input logic data_rvalid_i_1,
  input logic data_rvalid_i_2,
  input logic data_rvalidpar_i_1,
  input logic data_rvalidpar_i_2,
  output logic[31:0] data_wdata_o_1,
  output logic[31:0] data_wdata_o_2,
  output logic data_we_o_1,
  output logic data_we_o_2,
  output logic debug_halted_o_1,
  output logic debug_halted_o_2,
  output logic debug_havereset_o_1,
  output logic debug_havereset_o_2,
  output logic[31:0] debug_pc_o_1,
  output logic[31:0] debug_pc_o_2,
  output logic debug_pc_valid_o_1,
  output logic debug_pc_valid_o_2,
  input logic debug_req_i_1,
  input logic debug_req_i_2,
  output logic debug_running_o_1,
  output logic debug_running_o_2,
  input logic[31:0] dm_exception_addr_i_1,
  input logic[31:0] dm_exception_addr_i_2,
  input logic[31:0] dm_halt_addr_i_1,
  input logic[31:0] dm_halt_addr_i_2,
  input logic fencei_flush_ack_i_1,
  input logic fencei_flush_ack_i_2,
  output logic fencei_flush_req_o_1,
  output logic fencei_flush_req_o_2,
  input logic fetch_enable_i_1,
  input logic fetch_enable_i_2,
  output logic[12:0] instr_achk_o_1,
  output logic[12:0] instr_achk_o_2,
  output logic[31:0] instr_addr_o_1,
  output logic[31:0] instr_addr_o_2,
  output logic instr_dbg_o_1,
  output logic instr_dbg_o_2,
  input logic instr_err_i_1,
  input logic instr_err_i_2,
  input logic instr_gnt_i_1,
  input logic instr_gnt_i_2,
  input logic instr_gntpar_i_1,
  input logic instr_gntpar_i_2,
  output logic[1:0] instr_memtype_o_1,
  output logic[1:0] instr_memtype_o_2,
  output logic[2:0] instr_prot_o_1,
  output logic[2:0] instr_prot_o_2,
  input logic[4:0] instr_rchk_i_1,
  input logic[4:0] instr_rchk_i_2,
  input logic[31:0] instr_rdata_i_1,
  input logic[31:0] instr_rdata_i_2,
  output logic instr_req_o_1,
  output logic instr_req_o_2,
  output logic instr_reqpar_o_1,
  output logic instr_reqpar_o_2,
  input logic instr_rvalid_i_1,
  input logic instr_rvalid_i_2,
  input logic instr_rvalidpar_i_1,
  input logic instr_rvalidpar_i_2,
  input logic[31:0] irq_i_1,
  input logic[31:0] irq_i_2,
  output logic[63:0] mcycle_o_1,
  output logic[63:0] mcycle_o_2,
  input logic[31:0] mhartid_i_1,
  input logic[31:0] mhartid_i_2,
  input logic[3:0] mimpid_patch_i_1,
  input logic[3:0] mimpid_patch_i_2,
  input logic[31:0] mtvec_addr_i_1,
  input logic[31:0] mtvec_addr_i_2,
  input logic scan_cg_en_i_1,
  input logic scan_cg_en_i_2,
  input logic wu_wfe_i_1,
  input logic wu_wfe_i_2
);

logic rst_n;
assign rst_n = !rst;

cv32e40s_core U1(
  .alert_major_o(alert_major_o_1),
  .alert_minor_o(alert_minor_o_1),
  .boot_addr_i(boot_addr_i_1),
  .clic_irq_i(clic_irq_i_1),
  .clic_irq_id_i(clic_irq_id_i_1),
  .clic_irq_level_i(clic_irq_level_i_1),
  .clic_irq_priv_i(clic_irq_priv_i_1),
  .clic_irq_shv_i(clic_irq_shv_i_1),
  .clk_i(clk),
  .core_sleep_o(core_sleep_o_1),
  .data_achk_o(data_achk_o_1),
  .data_addr_o(data_addr_o_1),
  .data_be_o(data_be_o_1),
  .data_dbg_o(data_dbg_o_1),
  .data_err_i(data_err_i_1),
  .data_gnt_i(data_gnt_i_1),
  .data_gntpar_i(data_gntpar_i_1),
  .data_memtype_o(data_memtype_o_1),
  .data_prot_o(data_prot_o_1),
  .data_rchk_i(data_rchk_i_1),
  .data_rdata_i(data_rdata_i_1),
  .data_req_o(data_req_o_1),
  .data_reqpar_o(data_reqpar_o_1),
  .data_rvalid_i(data_rvalid_i_1),
  .data_rvalidpar_i(data_rvalidpar_i_1),
  .data_wdata_o(data_wdata_o_1),
  .data_we_o(data_we_o_1),
  .debug_halted_o(debug_halted_o_1),
  .debug_havereset_o(debug_havereset_o_1),
  .debug_pc_o(debug_pc_o_1),
  .debug_pc_valid_o(debug_pc_valid_o_1),
  .debug_req_i(debug_req_i_1),
  .debug_running_o(debug_running_o_1),
  .dm_exception_addr_i(dm_exception_addr_i_1),
  .dm_halt_addr_i(dm_halt_addr_i_1),
  .fencei_flush_ack_i(fencei_flush_ack_i_1),
  .fencei_flush_req_o(fencei_flush_req_o_1),
  .fetch_enable_i(fetch_enable_i_1),
  .instr_achk_o(instr_achk_o_1),
  .instr_addr_o(instr_addr_o_1),
  .instr_dbg_o(instr_dbg_o_1),
  .instr_err_i(instr_err_i_1),
  .instr_gnt_i(instr_gnt_i_1),
  .instr_gntpar_i(instr_gntpar_i_1),
  .instr_memtype_o(instr_memtype_o_1),
  .instr_prot_o(instr_prot_o_1),
  .instr_rchk_i(instr_rchk_i_1),
  .instr_rdata_i(instr_rdata_i_1),
  .instr_req_o(instr_req_o_1),
  .instr_reqpar_o(instr_reqpar_o_1),
  .instr_rvalid_i(instr_rvalid_i_1),
  .instr_rvalidpar_i(instr_rvalidpar_i_1),
  .irq_i(irq_i_1),
  .mcycle_o(mcycle_o_1),
  .mhartid_i(mhartid_i_1),
  .mimpid_patch_i(mimpid_patch_i_1),
  .mtvec_addr_i(mtvec_addr_i_1),
  .rst_ni(rst_n),
  .scan_cg_en_i(scan_cg_en_i_1),
  .wu_wfe_i(wu_wfe_i_1)
);

cv32e40s_core U2(
  .alert_major_o(alert_major_o_2),
  .alert_minor_o(alert_minor_o_2),
  .boot_addr_i(boot_addr_i_2),
  .clic_irq_i(clic_irq_i_2),
  .clic_irq_id_i(clic_irq_id_i_2),
  .clic_irq_level_i(clic_irq_level_i_2),
  .clic_irq_priv_i(clic_irq_priv_i_2),
  .clic_irq_shv_i(clic_irq_shv_i_2),
  .clk_i(clk),
  .core_sleep_o(core_sleep_o_2),
  .data_achk_o(data_achk_o_2),
  .data_addr_o(data_addr_o_2),
  .data_be_o(data_be_o_2),
  .data_dbg_o(data_dbg_o_2),
  .data_err_i(data_err_i_2),
  .data_gnt_i(data_gnt_i_2),
  .data_gntpar_i(data_gntpar_i_2),
  .data_memtype_o(data_memtype_o_2),
  .data_prot_o(data_prot_o_2),
  .data_rchk_i(data_rchk_i_2),
  .data_rdata_i(data_rdata_i_2),
  .data_req_o(data_req_o_2),
  .data_reqpar_o(data_reqpar_o_2),
  .data_rvalid_i(data_rvalid_i_2),
  .data_rvalidpar_i(data_rvalidpar_i_2),
  .data_wdata_o(data_wdata_o_2),
  .data_we_o(data_we_o_2),
  .debug_halted_o(debug_halted_o_2),
  .debug_havereset_o(debug_havereset_o_2),
  .debug_pc_o(debug_pc_o_2),
  .debug_pc_valid_o(debug_pc_valid_o_2),
  .debug_req_i(debug_req_i_2),
  .debug_running_o(debug_running_o_2),
  .dm_exception_addr_i(dm_exception_addr_i_2),
  .dm_halt_addr_i(dm_halt_addr_i_2),
  .fencei_flush_ack_i(fencei_flush_ack_i_2),
  .fencei_flush_req_o(fencei_flush_req_o_2),
  .fetch_enable_i(fetch_enable_i_2),
  .instr_achk_o(instr_achk_o_2),
  .instr_addr_o(instr_addr_o_2),
  .instr_dbg_o(instr_dbg_o_2),
  .instr_err_i(instr_err_i_2),
  .instr_gnt_i(instr_gnt_i_2),
  .instr_gntpar_i(instr_gntpar_i_2),
  .instr_memtype_o(instr_memtype_o_2),
  .instr_prot_o(instr_prot_o_2),
  .instr_rchk_i(instr_rchk_i_2),
  .instr_rdata_i(instr_rdata_i_2),
  .instr_req_o(instr_req_o_2),
  .instr_reqpar_o(instr_reqpar_o_2),
  .instr_rvalid_i(instr_rvalid_i_2),
  .instr_rvalidpar_i(instr_rvalidpar_i_2),
  .irq_i(irq_i_2),
  .mcycle_o(mcycle_o_2),
  .mhartid_i(mhartid_i_2),
  .mimpid_patch_i(mimpid_patch_i_2),
  .mtvec_addr_i(mtvec_addr_i_2),
  .rst_ni(rst_n),
  .scan_cg_en_i(scan_cg_en_i_2),
  .wu_wfe_i(wu_wfe_i_2)
);

endmodule // cv32e40s_miter
